*jk flip flop

.param Vdd=5  
Vdd Vdd 0 dc 5
MN1 1 clk 0 0 NCH L=0.18U     W=0.000.54996186000000
MN2 2 Q 1 0 NCH L=0.18U       W=0.000.19283916700000
MN3 3 K 2 0 NCH L=0.18U       W=0.000.1092328700000
MN4 4 3 0 0 NCH L=0.18U       W=0.000.65823972000000
MN5 O Q 4 0 NCH L=0.18U       W=0.00-0.9657540000000
MN6 6 clk 0 0 NCH L=0.18U     W=0.000.39184482000000
MN7 7 O 6 0 NCH L=0.18U       W=0.000.70053311400000
MN8 8 J 7 0 NCH L=0.18U       W=0.000.843967826000000
MP1 3 K Vdd Vdd PCH L=0.18U   W=0.000.976069802000000
MP2 3 Q Vdd Vdd PCH L=0.18U   W=0.00-0.2505029000000
MP3 3 clk Vdd Vdd PCH L=0.18U W=0.002.39518695000000
MP4 O 3  Vdd Vdd PCH L=0.18U  W=0.001.815404810000000
MP5 O Q Vdd Vdd PCH L=0.18U   W=0.00-0.034747770000
MP6 8 J Vdd Vdd PCH L=0.18U   W=0.000.705697301000000
MP7 8 O Vdd Vdd PCH L=0.18U   W=0.000.74332958000000
MP8 8 clk Vdd Vdd PCH L=0.18U W=0.000.520675570000000
MN9 17 8 0 0 NCH L=0.18U      W=0.001.25549613000000
MNN Q O 17 0 NCH L=0.18U      W=0.001.04419219400000
MP9 Q 8 Vdd Vdd PCH L=0.18U   W=0.000.0083942030000
MPP Q O Vdd Vdd PCH L=0.18U   W=0.000.226808439000

.MODEL PCH PMOS LEVEL=49
.MODEL NCH NMOS LEVEL=49

VJ J 0 PULSE 0 5 0 1N 1N 20N 40N
VK K 0 PULSE 0 5 20N 1N 1N 20N 40N
Vclk clk 0 PULSE 0 5 0 1N 1N 50N 100N

.MEASURE TRAN tplh TRIG V(j) VAL='Vdd/2' FALL=1 TARG V(Q)  VAL='Vdd/2'  FALL=1
.MEASURE TRAN tphl TRIG V(J) VAL='Vdd/2' RISE=2 TARG V(Q)  VAL='Vdd/2'  RISE=2
.MEASURE TRAN tPD PARAM='(tplh + tphl)/2'
.MEASURE TRAN tr TRIG V(Q) VAL='0.1*Vdd' RISE=1 TARG V(Q)  VAL='0.9*Vdd'  RISE=3
.MEASURE TRAN tf TRIG V(Q) VAL='0.9*Vdd' FALL=2 TARG V(Q)  VAL='0.1*Vdd'  FALL=1
.MEASURE TRAN tD PARAM='(tr + tf)/2' 

.meas tran AvgPower Avg Power from = 0ps to = 40ns
.meas tran maxpower max Power

.TRAN 1NS 200NS
.PRINT TRAN V(J) V(K) V(clk) V(Q) V(O)
.END